module mul (input [31:0] a,
		output [31:0] s) ;

assign s = 4 * a;

endmodule 